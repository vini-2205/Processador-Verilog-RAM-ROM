library verilog;
use verilog.vl_types.all;
entity test_pratica2 is
end test_pratica2;
